module inverter (output OUT, input IN);

	assign OUT = ~IN;

endmodule