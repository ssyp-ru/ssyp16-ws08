module not_16(input [15:0] A,output [15:0] RES);
assign RES=~A;
endmodule