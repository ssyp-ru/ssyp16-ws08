module cu();
	
endmodule
