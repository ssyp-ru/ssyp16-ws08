module part2()