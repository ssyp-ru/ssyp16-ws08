module memory (input [7:0] adress, output [15:0] op);


endmodule
