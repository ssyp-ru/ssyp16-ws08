module BC (input z, input [3:0] from_cu, input [3:0] from_fu, output [3:0] to_pc);


endmodule
