module multiplexor_offset(output [15:0] offset, input [15:0] imm_offset, input [15:0] A_offset)