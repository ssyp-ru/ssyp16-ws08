module and_16(input [15:0] A,input [15:0] B,output [15:0] RES);
assign RES=A & B;
endmodule