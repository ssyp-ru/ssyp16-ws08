//module main