module branch_control(output [15:0] N, input Z, input signal);
	always begin
		if (signal) begin
			
		end
	end
endmodule
