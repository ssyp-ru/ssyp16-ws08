module not_clk(output B, input A);
	assign B = ~A;
endmodule
