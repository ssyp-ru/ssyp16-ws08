module program_counter(output reg [7:0] pointer, input clk, input offset);

endmodule
